module Timer(
    reset_n, clk,
    timer_
);
endmodule