`timescale 1ns/1ns
`define PERIOD1 100
`define MEMORY_SIZE 256	//	size of memory is 2^8 words (reduced size)
`define WORD_SIZE 16	//	instead of 2^16 words to reduce memory
			//	requirements in the Active-HDL simulator 

module memory(clk, reset_n, read_m, write_m, address, data);
	input clk;
	wire clk;
	input reset_n;
	wire reset_n;
	
	input read_m;
	wire read_m;
	input write_m;
	wire write_m;
	input [`WORD_SIZE-1:0] address;
	wire [`WORD_SIZE-1:0] address;
	inout data;
	wire [`WORD_SIZE-1:0] data;
	
	reg [`WORD_SIZE-1:0] memory [0:`MEMORY_SIZE-1];
	reg [`WORD_SIZE-1:0] output_data;
	
	assign data = read_m?output_data:`WORD_SIZE'bz;
	
	always@(posedge clk)
		if(!reset_n)
			begin
				memory[16'h0] <= 16'h9023; // JMP
				memory[16'h1] <= 16'h1; // BNE
				memory[16'h2] <= 16'hffff; // R Type
				memory[16'h3] <= 16'h0; // BNE
				memory[16'h4] <= 16'h0; // BNE
				memory[16'h5] <= 16'h0; // BNE
				memory[16'h6] <= 16'h0; // BNE
				memory[16'h7] <= 16'h0; // BNE
				memory[16'h8] <= 16'h0; // BNE
				memory[16'h9] <= 16'h0; // BNE
				memory[16'ha] <= 16'h0; // BNE
				memory[16'hb] <= 16'h0; // BNE
				memory[16'hc] <= 16'h0; // BNE
				memory[16'hd] <= 16'h0; // BNE
				memory[16'he] <= 16'h0; // BNE
				memory[16'hf] <= 16'h0; // BNE
				memory[16'h10] <= 16'h0; // BNE
				memory[16'h11] <= 16'h0; // BNE
				memory[16'h12] <= 16'h0; // BNE
				memory[16'h13] <= 16'h0; // BNE
				memory[16'h14] <= 16'h0; // BNE
				memory[16'h15] <= 16'h0; // BNE
				memory[16'h16] <= 16'h0; // BNE
				memory[16'h17] <= 16'h0; // BNE
				memory[16'h18] <= 16'h0; // BNE
				memory[16'h19] <= 16'h0; // BNE
				memory[16'h1a] <= 16'h0; // BNE
				memory[16'h1b] <= 16'h0; // BNE
				memory[16'h1c] <= 16'h0; // BNE
				memory[16'h1d] <= 16'h0; // BNE
				memory[16'h1e] <= 16'h0; // BNE
				memory[16'h1f] <= 16'h0; // BNE
				memory[16'h20] <= 16'h0; // BNE
				memory[16'h21] <= 16'h0; // BNE
				memory[16'h22] <= 16'h0; // BNE
				memory[16'h23] <= 16'h6000;  // LHI 0
				memory[16'h24] <= 16'hf01c; // R Type
				memory[16'h25] <= 16'h6100; // LHI
				memory[16'h26] <= 16'hf41c; // R Type
				memory[16'h27] <= 16'h6200; // LHI
				memory[16'h28] <= 16'hf81c; // R Type
				memory[16'h29] <= 16'h6300; // LHI
				memory[16'h2a] <= 16'hfc1c; // R Type
				memory[16'h2b] <= 16'h4401; // 10. reg[0] = reg[1] + 1
				memory[16'h2c] <= 16'hf01c; // 11. WWD $0
				memory[16'h2d] <= 16'h4001; // ADI
				memory[16'h2e] <= 16'hf01c; // R Type
				memory[16'h2f] <= 16'h5901; // ODI
				memory[16'h30] <= 16'hf41c; // R Type
				memory[16'h31] <= 16'h5502; // ODI
				memory[16'h32] <= 16'hf41c; // R Type
				memory[16'h33] <= 16'h5503; // ODI
				memory[16'h34] <= 16'hf41c; // R Type
				memory[16'h35] <= 16'hf2c0; // R Type
				memory[16'h36] <= 16'hfc1c; // R Type
				memory[16'h37] <= 16'hf6c0; // R Type
				memory[16'h38] <= 16'hfc1c; // R Type
				memory[16'h39] <= 16'hf1c0; // R Type
				memory[16'h3a] <= 16'hfc1c; // R Type
				memory[16'h3b] <= 16'hf2c1; // R Type
				memory[16'h3c] <= 16'hfc1c; // R Type
				memory[16'h3d] <= 16'hf8c1; // R Type
				memory[16'h3e] <= 16'hfc1c; // R Type
				memory[16'h3f] <= 16'hf6c1; // R Type
				memory[16'h40] <= 16'hfc1c; // R Type
				memory[16'h41] <= 16'hf9c1; // R Type
				memory[16'h42] <= 16'hfc1c; // R Type
				memory[16'h43] <= 16'hf1c1; // R Type
				memory[16'h44] <= 16'hfc1c; // R Type
				memory[16'h45] <= 16'hf4c1; // R Type
				memory[16'h46] <= 16'hfc1c; // R Type
				memory[16'h47] <= 16'hf2c2; // R Type
				memory[16'h48] <= 16'hfc1c; // R Type
				memory[16'h49] <= 16'hf6c2; // R Type
				memory[16'h4a] <= 16'hfc1c; // R Type
				memory[16'h4b] <= 16'hf1c2; // R Type
				memory[16'h4c] <= 16'hfc1c; // R Type
				memory[16'h4d] <= 16'hf2c3; // R Type
				memory[16'h4e] <= 16'hfc1c; // R Type
				memory[16'h4f] <= 16'hf6c3; // R Type
				memory[16'h50] <= 16'hfc1c; // R Type
				memory[16'h51] <= 16'hf1c3; // R Type
				memory[16'h52] <= 16'hfc1c; // R Type
				memory[16'h53] <= 16'hf0c4; // R Type
				memory[16'h54] <= 16'hfc1c; // R Type
				memory[16'h55] <= 16'hf4c4; // R Type
				memory[16'h56] <= 16'hfc1c; // R Type
				memory[16'h57] <= 16'hf8c4; // R Type
				memory[16'h58] <= 16'hfc1c; // R Type
				memory[16'h59] <= 16'hf0c5; // R Type
				memory[16'h5a] <= 16'hfc1c; // R Type
				memory[16'h5b] <= 16'hf4c5; // R Type
				memory[16'h5c] <= 16'hfc1c; // R Type
				memory[16'h5d] <= 16'hf8c5; // R Type
				memory[16'h5e] <= 16'hfc1c; // R Type
				memory[16'h5f] <= 16'hf0c6; // R Type
				memory[16'h60] <= 16'hfc1c; // R Type
				memory[16'h61] <= 16'hf4c6; // R Type
				memory[16'h62] <= 16'hfc1c; // R Type
				memory[16'h63] <= 16'hf8c6; // R Type
				memory[16'h64] <= 16'hfc1c; // R Type
				memory[16'h65] <= 16'hf0c7; // R Type
				memory[16'h66] <= 16'hfc1c; // R Type
				memory[16'h67] <= 16'hf4c7; // R Type
				memory[16'h68] <= 16'hfc1c; // R Type
				memory[16'h69] <= 16'hf8c7; // R Type
				memory[16'h6a] <= 16'hfc1c; // R Type
				memory[16'h6b] <= 16'h7801; // LWD
				memory[16'h6c] <= 16'hf01c; // R Type
				memory[16'h6d] <= 16'h7902; // LWD
				memory[16'h6e] <= 16'hf41c; // R Type
				memory[16'h6f] <= 16'h8901; // SWD
				memory[16'h70] <= 16'h8802; // SWD
				memory[16'h71] <= 16'h7801; // LWD
				memory[16'h72] <= 16'hf01c; // R Type
				memory[16'h73] <= 16'h7902; // LWD
				memory[16'h74] <= 16'hf41c; // R Type
				memory[16'h75] <= 16'h9076; // JMP
				memory[16'h76] <= 16'hf01c; // R Type
				memory[16'h77] <= 16'h9079; // JMP
				memory[16'h78] <= 16'hf01d; // R Type
				memory[16'h79] <= 16'hf41c; // R Type
				memory[16'h7a] <= 16'hb01; // BNE
				memory[16'h7b] <= 16'h907d; // JMP
				memory[16'h7c] <= 16'hf01d; // R Type
				memory[16'h7d] <= 16'hf01c; // WWD 
				memory[16'h7e] <= 16'h601; // BNE
				memory[16'h7f] <= 16'hf01d; // R Type
				memory[16'h80] <= 16'hf41c; // R Type
				memory[16'h81] <= 16'h1601; // BEQ
				memory[16'h82] <= 16'h9084; // JMP
				memory[16'h83] <= 16'hf01d; // R Type
				memory[16'h84] <= 16'hf01c; // R Type
				memory[16'h85] <= 16'h1b01; // BEQ
				memory[16'h86] <= 16'hf01d; // R Type
				memory[16'h87] <= 16'hf41c; // R Type
				memory[16'h88] <= 16'h2001; // BGZ
				memory[16'h89] <= 16'h908b; // JMP
				memory[16'h8a] <= 16'hf01d; // R Type
				memory[16'h8b] <= 16'hf01c; // R Type
				memory[16'h8c] <= 16'h2401; // BGZ
				memory[16'h8d] <= 16'hf01d; // R Type
				memory[16'h8e] <= 16'hf41c; // R Type
				memory[16'h8f] <= 16'h2801; // BGZ
				memory[16'h90] <= 16'h9092; // JMP
				memory[16'h91] <= 16'hf01d; // R Type
				memory[16'h92] <= 16'hf01c; // R Type
				memory[16'h93] <= 16'h3001; // BLZ
				memory[16'h94] <= 16'hf01d; // R Type
				memory[16'h95] <= 16'hf41c; // R Type
				memory[16'h96] <= 16'h3401; // BLZ
				memory[16'h97] <= 16'h9099; // JMP
				memory[16'h98] <= 16'hf01d; // R Type
				memory[16'h99] <= 16'hf01c; // R Type
				memory[16'h9a] <= 16'h3801; // BLZ
				memory[16'h9b] <= 16'h909d; // JMP
				memory[16'h9c] <= 16'hf01d; // R Type
				memory[16'h9d] <= 16'hf41c; // R Type WWD
				memory[16'h9e] <= 16'ha0af; // JAL ****************
				memory[16'h9f] <= 16'hf01c; // R Type
				memory[16'ha0] <= 16'ha0ae; // JAL
				memory[16'ha1] <= 16'hf01d; // R Type
				memory[16'ha2] <= 16'hf41c; // R Type
				memory[16'ha3] <= 16'h6300; // LHI
				memory[16'ha4] <= 16'h5f03; // ODI
				memory[16'ha5] <= 16'h6000; // LHI
				memory[16'ha6] <= 16'h4005; // ADI
				memory[16'ha7] <= 16'ha0b2; // JAL
				memory[16'ha8] <= 16'hf01c; // R Type
				memory[16'ha9] <= 16'h90b1; // JMP
				memory[16'haa] <= 16'h4900; // ADI
				memory[16'hab] <= 16'hf41a; // R Type
				memory[16'hac] <= 16'hf01c; // R Type
				memory[16'had] <= 16'hf01d; // R Type
				memory[16'hae] <= 16'h4a01; // ADI
				memory[16'haf] <= 16'hf819; // R Type
				memory[16'hb0] <= 16'hf01d; // R Type
				memory[16'hb1] <= 16'ha0aa; // JAL
				memory[16'hb2] <= 16'h41ff; // ADI
				memory[16'hb3] <= 16'h2404; // BGZ
				memory[16'hb4] <= 16'h6000; // LHI
				memory[16'hb5] <= 16'h5001; // ODI
				memory[16'hb6] <= 16'hf819; // R Type
				memory[16'hb7] <= 16'hf01d; // R Type
				memory[16'hb8] <= 16'h8e00; // SWD
				memory[16'hb9] <= 16'h8c01; // SWD
				memory[16'hba] <= 16'h4f02; // ADI
				memory[16'hbb] <= 16'h40fe; // ADI
				memory[16'hbc] <= 16'ha0b2; // JAL
				memory[16'hbd] <= 16'h7dff; // LWD
				memory[16'hbe] <= 16'h8cff; // SWD
				memory[16'hbf] <= 16'h44ff; // ADI
				memory[16'hc0] <= 16'ha0b2; // JAL
				memory[16'hc1] <= 16'h7dff; // LWD
				memory[16'hc2] <= 16'h7efe; // LWD
				memory[16'hc3] <= 16'hf100; // R Type
				memory[16'hc4] <= 16'h4ffe; // ADI
				memory[16'hc5] <= 16'hf819; // R Type
				memory[16'hc6] <= 16'hf01d; // R Type
			end
		else
			begin
				if(read_m)output_data <= memory[address];
				if(write_m)memory[address] <= data;
			end
endmodule